`include "gsf.svh"

module hw_top;

integer id = 0;

`gsf_is_buf(DataQ, 512,12);

endmodule
